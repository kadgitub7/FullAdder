`timescale 1ns / 1ps

module fulladder(
    input A,
    input B,
    input Ci,
    output S,
    output Co
    );
    
    assign S = A^B^Ci;
    assign Co = A&B | A&Ci | B&Ci;
endmodule